module ALU #(parameter bus_size) (input logic[bus_size-1:0] a, b, input logic[2:0]c, 
											output logic[bus_size-1:0] s, output logic flag_overflow, flag_zero, 
											flag_negative, flag_carry);
	
		
		
endmodule
